`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   17:29:26 03/28/2007
// Design Name:   f1
// Module Name:   test.v
// Project Name:  sudokuf1
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: f1
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module test_v;

	// Inputs
	reg clock;
	reg [1:810] arri;
	reg load;

	// Outputs
	wire done;
	wire [1:810] arro;
	integer i;
//	wire [1:81] temp1, temp2, temp3;
//	wire [1:729] temp;
//	wire [1:729] ftemp1, ftemp2, ftemp3, f1temp, f2temp2, f2temp;
	

	// Instantiate the Unit Under Test (UUT)
	f1 uut (
		.clock(clock), 
		.arri(arri), 
		.done(done), 
		.load(load), 
		.arro(arro)
	//	.temp1(temp1),
	//	.temp2(temp2),
	//	.temp3(temp3),
	//	.f1temp(f1temp), 
	//	.ftemp1(ftemp1), 
	//	.ftemp2(ftemp2), 
	//	.ftemp3(ftemp3), 
	//	.f2temp2(f2temp2), 
	//	.f2temp(f2temp),
	//	.temp(temp)
	);

	initial begin
		// Initialize Inputs
		clock = 0;
		arri = 0;
		load = 0;

		 $dumpfile("sudokuf1.vcd"); // save waveforms in this file
     $dumpvars;  // saves all waveforms


	#2 load = 1;
	
	//first: 8 Cycles
//	#2 arri = 810'b000000000010000000010000000000000000000000000000000000010001000100000101000000010000000101000000000000000000000000000000000010000100000000000010000001000000000000000000000000010001000000000000000100010001000001010000000100000000000000000000001000000100000000000000100001100000000100000010010000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000100001000000000000000001010000000000010000000100000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000010011000000001001000000100000000001000000001000000000000000000000100000001000001000100000001010000000000000000010100000000000000000000000000100100000000001000000001000000000000000000000000000000000100000101000000010000001001000000010100000000000000000000000000000000001000010000000000;
	//fourth: 12 cycles
//	#2 arri = 810'b000000000000000000000000000011000010000100000000000000000000000100000100000000000000000000000000000010000000010000000000000000000000000000000000000000000000001100000001010000000000000000000000010000010000100001000000000000000001010000000000001000000100000000000100000001000000000000000000001000000001001000000100000000000000010001000000000000000000000000000000000000000000000010010000000000000000010100000000110000100001000000000001000000010000000000000000000000000000000000000000000000100100000000000001000001000010000100000000000000000000010000000100000000000000000101000000000000010000010000000000000001000100001000010000000000000000000000001000010001000001000000000000000000000000000000000000000000000000110000000000000000000000000000000000001001000000000000000000000010000001010000000100000000000000000000;
	//final: 11 cycles
//	#2 arri = 810'b000000100100000001010000000000000000000000000000000000100001000000000000100000010001000001000000000000000000000000000000000000000000000000000000000000000010000100000010010000000000000000000000000000000000000000001000000100000000000000000000000000001101000000010000000000000010000110000000010000000011000000000000000000000000001001000000000000000000000000000000000001000100000000000000000000000000000000000000000000000000000000000000000000000000000011000000000000000000000000000000000100000100000000000000000000100000000100001000010100000001000000000000001000010100000001000000000000000000001000000001000000000000000000000000000000000000000000010000010000010001000000000000000000000000000000000000000000000000000000000000100000000100000010010000000000000000001100000000000000000000000000000000000100010000100001;		
	//second: 10 cycles
//	#2 arri = 810'b000000100100000000000000000000000000000000000100010000000000010000000100100000010000000000000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000001010000100001010000000110000000010000000000000100000100000100010000000000000000001100000010011000000001000000000000001000010000010001000000000000000000000000000000000000000000010000010000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000100000000100000000110000000000000001000100010000010000001001000000000000001000010000001001000000000000000001010000000011001000000110000000010000000000000000000000000000000000000000000000000001000000010000000000000000000000000000000000000000000000000010000000010000000011000000000000000010010000000000000000000000000000000100000001;
	//third: 7 cycles
	#2 arri = 810'b000000000000000000000000000000001000000100000000000000000000100000000100000000110000000000000000000000000000000000000011000000000000000010010000000000000000010100000000000000010001000000000000000000001000000001000000000000000100010000000000000000000000001000010100000001001000000100000001010000000000010000000100000000110000000000000000000000000000000000000000000000000000000010010000100001000001000100000000000000000101010000000100100000010000000000000000000000000000000000000000000000000000100000011000000001000000000000000001010000100001000000001100001000010000000000000000000010000000010000000000000001000100000000000000000000010000000100000000000000001001000000000000000001010000000000000010000100000000000000000000000000000010000000010010000001000000000000000000000000010001000000000000000000000000000000;
	
	#12 load = 0;	

#200 for (i=1; i<=810; i=i+1)
     begin
     	$write(arro[i]);
	if ((i%10) == 0)
		$write(" ");
	if ((i%90) == 0)
		$write("\n");
     end

#2 $finish;
	end
	
	always #2 clock = ~clock;
      
endmodule



