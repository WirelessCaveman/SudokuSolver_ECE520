module f1 (clock, arri, done, load, arro/*, temp1, temp2, temp3, f1temp, ftemp1,
ftemp2, ftemp3, f2temp2, f2temp, temp*/);
	input clock; // Clock
	input [1:810] arri;
	input load;
	
	// all outputs are registered
	output done;
	output [1:810] arro;
//	output [1:81] temp1, temp2, temp3;
//	output [1:729] temp; 
//	output [1:729] ftemp1, ftemp2, ftemp3, f1temp, f2temp, f2temp2;
	
	integer i, j, x;
	reg [1:81] temp1, temp2, temp3;
	reg [1:729] temp, f1temp, f2temp, f2temp2;
	reg [1:729] ftemp1, ftemp2, ftemp3;
	reg [1:810]arr;
	reg done;
	reg [1:810] arro;
	wire [1:810] arri;
	reg  count;
	
	always @ (posedge clock)
	begin
		if (load == 1)
		begin
			count <= 0;
		end
		else
		begin
			count <= ~(count);

		end
	end
	
	always@ (arr)	//for row
	begin
		for (i = 1; i < 10; i=i+1)
		begin
			for (x = 1; x < 10; x=x+1) //bit positions for same cell
			begin	
				temp1[(i-1)*9 + x] = |{(arr[(i-1)*90 + 0*10 + x] && arr[(i-1)*90 + 0*10 + 10]), (arr[(i-1)*90 + 1*10 + x] && arr[(i-1)*90 + 1*10 + 10]), (arr[(i-1)*90 + 2*10 + x] && arr[(i-1)*90 + 2*10 + 10]), (arr[(i-1)*90 + 3*10 + x] && arr[(i-1)*90 + 3*10 + 10]), (arr[(i-1)*90 + 4*10 + x] && arr[(i-1)*90 + 4*10 + 10]), (arr[(i-1)*90 + 5*10 + x] && arr[(i-1)*90 + 5*10 + 10]), (arr[(i-1)*90 + 6*10 + x] && arr[(i-1)*90 + 6*10 + 10]), (arr[(i-1)*90 + 7*10 + x] && arr[(i-1)*90 + 7*10 + 10]), (arr[(i-1)*90 + 8*10 + x] && arr[(i-1)*90 + 8*10 + 10])};
			end
		end
	end
	
	always @ (arr)	//for column
	begin
		for (i = 1; i < 10; i=i+1)
		begin
			for (x = 1; x < 10; x=x+1) //bit positions for same cell
			begin
				temp2[(i-1)*9 + x] = |{(arr[0*90 + (i-1)*10 + x] && arr[0*90 + (i-1)*10 + 10]), (arr[1*90 + (i-1)*10 + x] && arr[1*90 + (i-1)*10 + 10]), (arr[2*90 + (i-1)*10 + x] && arr[2*90 + (i-1)*10 + 10]), (arr[3*90 + (i-1)*10 + x] && arr[3*90 + (i-1)*10 + 10]), (arr[4*90 + (i-1)*10 + x] && arr[4*90 + (i-1)*10 + 10]), (arr[5*90 + (i-1)*10 + x] && arr[5*90 + (i-1)*10 + 10]), (arr[6*90 + (i-1)*10 + x] && arr[6*90 + (i-1)*10 + 10]), (arr[7*90 + (i-1)*10 + x] && arr[7*90 + (i-1)*10 + 10]), (arr[8*90 + (i-1)*10 + x] && arr[8*90 + (i-1)*10 + 10])};
			end
		end
	end
	
	always @ (arr)	//for square
	begin				
		for (i = 1; i < 10; i=i+1)
		begin	
			for (x = 1; x < 10; x = x+1)
			begin
				temp3[(i-1)*9 + x]= |{(arr[((i-1)/3)*270 + ((i-1)%3)*30 + 0 + x] && arr[((i-1)/3)*270 + ((i-1)%3)*30 + 0 + 10]), (arr[((i-1)/3)*270 + ((i-1)%3)*30 + 10 + x] && arr[((i-1)/3)*270 + ((i-1)%3)*30 + 10 + 10]), (arr[((i-1)/3)*270 + ((i-1)%3)*30 + 20 + x] && arr[((i-1)/3)*270 + ((i-1)%3)*30 + 20 + 10]),
									  (arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 0 + x] && arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 0 + 10]), (arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 10 + x] && arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 10 + 10]), (arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 20 + x] && arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 20 + 10]),
									  (arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + x] && arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + 10]), (arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 10 + x] && arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 10 + 10]), (arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 20 + x] && arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 20 + 10])};
			end
		end
	end	//always @
	
	always @ (temp1 or temp2 or temp3 or arr)	//combining row, column and square
	begin	
		for (i = 1; i < 82; i=i+1)
		begin
	 		if (arr[(i-1)*10 + 10] == 0)	//mux1: modified value from the combination logic to be selected- this cell is yet to be confirmed
			begin
	 			for (x = 1; x < 10; x=x+1) //bit positions for same cell
				begin
					f1temp[(i-1)*9 + x] = ~(|{temp1[((i-1)/9)*9 + x], temp2[((i-1)%9)*9 + x], temp3[(((i-1)/27)*3 + ((i-1)%9)/3)*9 + x]});
				end
			end
			else	//mux1: old value from the register should be selected since this cell is already confirmed
			begin
				for (x = 1; x < 10; x=x+1) 
				begin
					f1temp[(i-1)*9 + x] = arr[(i-1)*10 + x];
				end
			end
		end
	end	//always@		
		
		
	always @ (arr)
	begin
		for (i = 1; i < 82; i = i+1)
		begin
			for (x = 1; x < 11; x = x+1)
			begin
				arro[(i-1)*10 + x] = arr[(i-1)*10 + x];
			end
		end
		done = &{arr[(8*9 + 1)*10], arr[(8*9 + 2)*10], arr[(8*9 + 3)*10], arr[(8*9 + 4)*10], arr[(8*9 + 5)*10], arr[(8*9 + 6)*10], arr[(8*9 + 7)*10], arr[(8*9 + 8)*10], arr[(8*9 + 9)*10], 
				 arr[(7*9 + 1)*10], arr[(7*9 + 2)*10], arr[(7*9 + 3)*10], arr[(7*9 + 4)*10], arr[(7*9 + 5)*10], arr[(7*9 + 6)*10], arr[(7*9 + 7)*10], arr[(7*9 + 8)*10], arr[(7*9 + 9)*10], 
				 arr[(6*9 + 1)*10], arr[(6*9 + 2)*10], arr[(6*9 + 3)*10], arr[(6*9 + 4)*10], arr[(6*9 + 5)*10], arr[(6*9 + 6)*10], arr[(6*9 + 7)*10], arr[(6*9 + 8)*10], arr[(6*9 + 9)*10],
				 arr[(5*9 + 1)*10], arr[(5*9 + 2)*10], arr[(5*9 + 3)*10], arr[(5*9 + 4)*10], arr[(5*9 + 5)*10], arr[(5*9 + 6)*10], arr[(5*9 + 7)*10], arr[(5*9 + 8)*10], arr[(5*9 + 9)*10], 
				 arr[(4*9 + 1)*10], arr[(4*9 + 2)*10], arr[(4*9 + 3)*10], arr[(4*9 + 4)*10], arr[(4*9 + 5)*10], arr[(4*9 + 6)*10], arr[(4*9 + 7)*10], arr[(4*9 + 8)*10], arr[(4*9 + 9)*10], 
				 arr[(3*9 + 1)*10], arr[(3*9 + 2)*10], arr[(3*9 + 3)*10], arr[(3*9 + 4)*10], arr[(3*9 + 5)*10], arr[(3*9 + 6)*10], arr[(3*9 + 7)*10], arr[(3*9 + 8)*10], arr[(3*9 + 9)*10], 
				 arr[(2*9 + 1)*10], arr[(2*9 + 2)*10], arr[(2*9 + 3)*10], arr[(2*9 + 4)*10], arr[(2*9 + 5)*10], arr[(2*9 + 6)*10], arr[(2*9 + 7)*10], arr[(2*9 + 8)*10], arr[(2*9 + 9)*10], 
				 arr[(1*9 + 1)*10], arr[(1*9 + 2)*10], arr[(1*9 + 3)*10], arr[(1*9 + 4)*10], arr[(1*9 + 5)*10], arr[(1*9 + 6)*10], arr[(1*9 + 7)*10], arr[(1*9 + 8)*10], arr[(1*9 + 9)*10],
				 arr[(0*9 + 1)*10], arr[(0*9 + 2)*10], arr[(0*9 + 3)*10], arr[(0*9 + 4)*10], arr[(0*9 + 5)*10], arr[(0*9 + 6)*10], arr[(0*9 + 7)*10], arr[(0*9 + 8)*10], arr[(0*9 + 9)*10]};
	end
	
/******************************************************************************************/	
/*******************************            F2              *******************************/
/******************************************************************************************/

	always @ (arr)
	begin
		//for each row
		for (i = 1; i < 10; i=i+1)	//each i represents one row
		begin
			for (x = 1; x < 10; x=x+1)	//each x represents a bit position
			begin	
				ftemp1[(i-1)*81 + 0*9 + x] = (arr[(i-1)*90 + 0*10 + x] && (~|{arr[(i-1)*90 + 1*10 + x], arr[(i-1)*90 + 2*10 + x], arr[(i-1)*90 + 3*10 + x], arr[(i-1)*90 + 4*10 + x], arr[(i-1)*90 + 5*10 + x], arr[(i-1)*90 + 6*10 + x], arr[(i-1)*90 + 7*10 + x], arr[(i-1)*90 + 8*10 + x]})); 	//first cell in the row			[(i-1)*90 + x]
				ftemp1[(i-1)*81 + 1*9 + x] = (arr[(i-1)*90 + 1*10 + x] && (~|{arr[(i-1)*90 + 0*10 + x], arr[(i-1)*90 + 2*10 + x], arr[(i-1)*90 + 3*10 + x], arr[(i-1)*90 + 4*10 + x], arr[(i-1)*90 + 5*10 + x], arr[(i-1)*90 + 6*10 + x], arr[(i-1)*90 + 7*10 + x], arr[(i-1)*90 + 8*10 + x]})); 	//second cell in the row
				ftemp1[(i-1)*81 + 2*9 + x] = (arr[(i-1)*90 + 2*10 + x] && (~|{arr[(i-1)*90 + 0*10 + x], arr[(i-1)*90 + 1*10 + x], arr[(i-1)*90 + 3*10 + x], arr[(i-1)*90 + 4*10 + x], arr[(i-1)*90 + 5*10 + x], arr[(i-1)*90 + 6*10 + x], arr[(i-1)*90 + 7*10 + x], arr[(i-1)*90 + 8*10 + x]})); 	//third cell in the row
				ftemp1[(i-1)*81 + 3*9 + x] = (arr[(i-1)*90 + 3*10 + x] && (~|{arr[(i-1)*90 + 0*10 + x], arr[(i-1)*90 + 1*10 + x], arr[(i-1)*90 + 2*10 + x], arr[(i-1)*90 + 4*10 + x], arr[(i-1)*90 + 5*10 + x], arr[(i-1)*90 + 6*10 + x], arr[(i-1)*90 + 7*10 + x], arr[(i-1)*90 + 8*10 + x]})); 	//fourth cell in the row
				ftemp1[(i-1)*81 + 4*9 + x] = (arr[(i-1)*90 + 4*10 + x] && (~|{arr[(i-1)*90 + 0*10 + x], arr[(i-1)*90 + 1*10 + x], arr[(i-1)*90 + 2*10 + x], arr[(i-1)*90 + 3*10 + x], arr[(i-1)*90 + 5*10 + x], arr[(i-1)*90 + 6*10 + x], arr[(i-1)*90 + 7*10 + x], arr[(i-1)*90 + 8*10 + x]})); 	//fifth cell in the row
				ftemp1[(i-1)*81 + 5*9 + x] = (arr[(i-1)*90 + 5*10 + x] && (~|{arr[(i-1)*90 + 0*10 + x], arr[(i-1)*90 + 1*10 + x], arr[(i-1)*90 + 2*10 + x], arr[(i-1)*90 + 3*10 + x], arr[(i-1)*90 + 4*10 + x], arr[(i-1)*90 + 6*10 + x], arr[(i-1)*90 + 7*10 + x], arr[(i-1)*90 + 8*10 + x]})); 	//sixth cell in the row
				ftemp1[(i-1)*81 + 6*9 + x] = (arr[(i-1)*90 + 6*10 + x] && (~|{arr[(i-1)*90 + 0*10 + x], arr[(i-1)*90 + 1*10 + x], arr[(i-1)*90 + 2*10 + x], arr[(i-1)*90 + 3*10 + x], arr[(i-1)*90 + 4*10 + x], arr[(i-1)*90 + 5*10 + x], arr[(i-1)*90 + 7*10 + x], arr[(i-1)*90 + 8*10 + x]})); 	//seventh cell in the row
				ftemp1[(i-1)*81 + 7*9 + x] = (arr[(i-1)*90 + 7*10 + x] && (~|{arr[(i-1)*90 + 0*10 + x], arr[(i-1)*90 + 1*10 + x], arr[(i-1)*90 + 2*10 + x], arr[(i-1)*90 + 3*10 + x], arr[(i-1)*90 + 4*10 + x], arr[(i-1)*90 + 5*10 + x], arr[(i-1)*90 + 6*10 + x], arr[(i-1)*90 + 8*10 + x]})); 	//eighth cell in the row
				ftemp1[(i-1)*81 + 8*9 + x] = (arr[(i-1)*90 + 8*10 + x] && (~|{arr[(i-1)*90 + 0*10 + x], arr[(i-1)*90 + 1*10 + x], arr[(i-1)*90 + 2*10 + x], arr[(i-1)*90 + 3*10 + x], arr[(i-1)*90 + 4*10 + x], arr[(i-1)*90 + 5*10 + x], arr[(i-1)*90 + 6*10 + x], arr[(i-1)*90 + 7*10 + x]})); 	//ninth cell in the row
			end
		end
	end
	
	always @ (arr)
	begin
		//for each column
		for (i = 1; i < 10; i=i+1)	//each i represents one column
		begin
			for (x = 1; x < 10; x=x+1)	//each x represents a bit position
			begin	
				ftemp2[0*81 + (i-1)*9 + x] = (arr[0*90 + (i-1)*10 + x] && (~|{arr[(i-1)*10 + 1*90 + x], arr[(i-1)*10 + 2*90 + x], arr[(i-1)*10 + 3*90 + x], arr[(i-1)*10 + 4*90 + x], arr[(i-1)*10 + 5*90 + x], arr[(i-1)*10 + 6*90 + x], arr[(i-1)*10 + 7*90 + x], arr[(i-1)*10 + 8*90 + x]})); 	//first cell in the row			[(i-1)*10 + x]
				ftemp2[1*81 + (i-1)*9 + x] = (arr[1*90 + (i-1)*10 + x] && (~|{arr[(i-1)*10 + 0*90 + x], arr[(i-1)*10 + 2*90 + x], arr[(i-1)*10 + 3*90 + x], arr[(i-1)*10 + 4*90 + x], arr[(i-1)*10 + 5*90 + x], arr[(i-1)*10 + 6*90 + x], arr[(i-1)*10 + 7*90 + x], arr[(i-1)*10 + 8*90 + x]})); 	//second cell in the row
				ftemp2[2*81 + (i-1)*9 + x] = (arr[2*90 + (i-1)*10 + x] && (~|{arr[(i-1)*10 + 0*90 + x], arr[(i-1)*10 + 1*90 + x], arr[(i-1)*10 + 3*90 + x], arr[(i-1)*10 + 4*90 + x], arr[(i-1)*10 + 5*90 + x], arr[(i-1)*10 + 6*90 + x], arr[(i-1)*10 + 7*90 + x], arr[(i-1)*10 + 8*90 + x]})); 	//third cell in the row
				ftemp2[3*81 + (i-1)*9 + x] = (arr[3*90 + (i-1)*10 + x] && (~|{arr[(i-1)*10 + 0*90 + x], arr[(i-1)*10 + 1*90 + x], arr[(i-1)*10 + 2*90 + x], arr[(i-1)*10 + 4*90 + x], arr[(i-1)*10 + 5*90 + x], arr[(i-1)*10 + 6*90 + x], arr[(i-1)*10 + 7*90 + x], arr[(i-1)*10 + 8*90 + x]})); 	//fourth cell in the row
				ftemp2[4*81 + (i-1)*9 + x] = (arr[4*90 + (i-1)*10 + x] && (~|{arr[(i-1)*10 + 0*90 + x], arr[(i-1)*10 + 1*90 + x], arr[(i-1)*10 + 2*90 + x], arr[(i-1)*10 + 3*90 + x], arr[(i-1)*10 + 5*90 + x], arr[(i-1)*10 + 6*90 + x], arr[(i-1)*10 + 7*90 + x], arr[(i-1)*10 + 8*90 + x]})); 	//fifth cell in the row
				ftemp2[5*81 + (i-1)*9 + x] = (arr[5*90 + (i-1)*10 + x] && (~|{arr[(i-1)*10 + 0*90 + x], arr[(i-1)*10 + 1*90 + x], arr[(i-1)*10 + 2*90 + x], arr[(i-1)*10 + 3*90 + x], arr[(i-1)*10 + 4*90 + x], arr[(i-1)*10 + 6*90 + x], arr[(i-1)*10 + 7*90 + x], arr[(i-1)*10 + 8*90 + x]})); 	//sixth cell in the row
				ftemp2[6*81 + (i-1)*9 + x] = (arr[6*90 + (i-1)*10 + x] && (~|{arr[(i-1)*10 + 0*90 + x], arr[(i-1)*10 + 1*90 + x], arr[(i-1)*10 + 2*90 + x], arr[(i-1)*10 + 3*90 + x], arr[(i-1)*10 + 4*90 + x], arr[(i-1)*10 + 5*90 + x], arr[(i-1)*10 + 7*90 + x], arr[(i-1)*10 + 8*90 + x]})); 	//seventh cell in the row
				ftemp2[7*81 + (i-1)*9 + x] = (arr[7*90 + (i-1)*10 + x] && (~|{arr[(i-1)*10 + 0*90 + x], arr[(i-1)*10 + 1*90 + x], arr[(i-1)*10 + 2*90 + x], arr[(i-1)*10 + 3*90 + x], arr[(i-1)*10 + 4*90 + x], arr[(i-1)*10 + 5*90 + x], arr[(i-1)*10 + 6*90 + x], arr[(i-1)*10 + 8*90 + x]})); 	//eighth cell in the row
				ftemp2[8*81 + (i-1)*9 + x] = (arr[8*90 + (i-1)*10 + x] && (~|{arr[(i-1)*10 + 0*90 + x], arr[(i-1)*10 + 1*90 + x], arr[(i-1)*10 + 2*90 + x], arr[(i-1)*10 + 3*90 + x], arr[(i-1)*10 + 4*90 + x], arr[(i-1)*10 + 5*90 + x], arr[(i-1)*10 + 6*90 + x], arr[(i-1)*10 + 7*90 + x]})); 	//ninth cell in the row
			end
		end
	end
	
	always @ (arr)
	begin
		//for each square
		for (i = 1; i < 10; i=i+1)	//each i represents one square
		begin
			for (x = 1; x < 10; x=x+1)	//each x represents a bit position
			begin
				ftemp3[((i-1)/3)*243 + ((i-1)%3)*27 + 0 + x]  = (arr[((i-1)/3)*270 + ((i-1)%3)*30 + 0 + x] && (~|{arr[((i-1)/3)*270 + ((i-1)%3)*30 + 10 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 20 + x]}));
				ftemp3[((i-1)/3)*243 + ((i-1)%3)*27 + 9 + x] = (arr[((i-1)/3)*270 + ((i-1)%3)*30 + 10 + x] && (~|{arr[((i-1)/3)*270 + ((i-1)%3)*30 + 0 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 20 + x]}));
				ftemp3[((i-1)/3)*243 + ((i-1)%3)*27 + 18 + x] = (arr[((i-1)/3)*270 + ((i-1)%3)*30 + 20 + x] && (~|{arr[((i-1)/3)*270 + ((i-1)%3)*30 + 0 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 20 + x]}));
				ftemp3[(((i-1)/3)*243) + 81 + ((i-1)%3)*27 + 0 + x]  = (arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 0 + x] && (~|{arr[((i-1)/3)*270 + ((i-1)%3)*30 + 0 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 10 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 20 + x]}));
				ftemp3[(((i-1)/3)*243) + 81 + ((i-1)%3)*27 + 9 + x] = (arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 10 + x] && (~|{arr[((i-1)/3)*270 + ((i-1)%3)*30 + 0 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 10 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 20 + x]}));
				ftemp3[(((i-1)/3)*243) + 81 + ((i-1)%3)*27 + 18 + x] = (arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 20 + x] && (~|{arr[((i-1)/3)*270 + ((i-1)%3)*30 + 0 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 10 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 20 + x]}));
				ftemp3[(((i-1)/3)*243) + 162 + ((i-1)%3)*27 + 0 + x] =  (arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + x] && (~|{arr[((i-1)/3)*270 + ((i-1)%3)*30 + 0 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 10 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 20 + x]}));
				ftemp3[(((i-1)/3)*243) + 162 + ((i-1)%3)*27 + 9 + x] = (arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + x] && (~|{arr[((i-1)/3)*270 + ((i-1)%3)*30 + 0 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 10 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 20 + x]}));
				ftemp3[(((i-1)/3)*243) + 162 + ((i-1)%3)*27 + 18 + x] = (arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + x] && (~|{arr[((i-1)/3)*270 + ((i-1)%3)*30 + 0 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 10 + x], arr[((i-1)/3)*270 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 10 + x], arr[(((i-1)/3)*270) + 90 + ((i-1)%3)*30 + 20 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 0 + x], arr[(((i-1)/3)*270) + 180 + ((i-1)%3)*30 + 10 + x]}));
			end
		end
	end
	
	always @ (ftemp1 or ftemp2 or ftemp3)
	begin
		for (i = 1; i < 730; i=i+1)
		begin
			f2temp2[i] = |{ftemp1[i], ftemp2[i], ftemp3[i]};
		end
	end
	
	always @ (f2temp2 or arr)
	begin
		for (i = 1; i < 82; i=i+1)
		begin
			if ({f2temp2[(i-1)*9 + 1], f2temp2[(i-1)*9 + 2], f2temp2[(i-1)*9 + 3], f2temp2[(i-1)*9 + 4], f2temp2[(i-1)*9 + 5], f2temp2[(i-1)*9 + 6], f2temp2[(i-1)*9 + 7], f2temp2[(i-1)*9 + 8], f2temp2[((i-1)*9 + 9)]} == 9'b0)
			begin
				{f2temp[(i-1)*9 + 1], f2temp[(i-1)*9 + 2], f2temp[(i-1)*9 + 3], f2temp[(i-1)*9 + 4], f2temp[(i-1)*9 + 5], f2temp[(i-1)*9 + 6], f2temp[(i-1)*9 + 7], f2temp[(i-1)*9 + 8], f2temp[((i-1)*9 + 9)]} = {arr[(i-1)*10 + 1], arr[(i-1)*10 + 2], arr[(i-1)*10 + 3], arr[(i-1)*10 + 4], arr[(i-1)*10 + 5], arr[(i-1)*10 + 6], arr[(i-1)*10 + 7], arr[(i-1)*10 + 8], arr[((i-1)*10 + 9)]};
			end
			else
			begin
				{f2temp[(i-1)*9 + 1], f2temp[(i-1)*9 + 2], f2temp[(i-1)*9 + 3], f2temp[(i-1)*9 + 4], f2temp[(i-1)*9 + 5], f2temp[(i-1)*9 + 6], f2temp[(i-1)*9 + 7], f2temp[(i-1)*9 + 8], f2temp[((i-1)*9 + 9)]} = {f2temp2[(i-1)*9 + 1], f2temp2[(i-1)*9 + 2], f2temp2[(i-1)*9 + 3], f2temp2[(i-1)*9 + 4], f2temp2[(i-1)*9 + 5], f2temp2[(i-1)*9 + 6], f2temp2[(i-1)*9 + 7], f2temp2[(i-1)*9 + 8], f2temp2[((i-1)*9 + 9)]};
			end
		end
	end
	
	
	/************************************************************************/
	/****************COMBINE F1 AND F2***************************************/
	/************************************************************************/
	
	always @ (count or f1temp or f2temp)
	begin
		if (count == 0)
		begin
			for (i = 1; i < 730; i=i+1)
			begin
				temp[i] = f1temp[i];
			end
		end
		else
		begin
			for (i = 1; i < 730; i=i+1)
			begin
				temp[i] =  f2temp[i];
			end
		end
	end
	
	always @ (posedge clock)
	begin		
			for (i = 1; i < 82; i = i+1)
			begin
				if (load == 1)	//mux2: load initial input values
				begin	
					for (x = 1; x < 11; x = x+1)
					begin
						arr[(i-1)*10 + x] <= arri[(i-1)*10 + x];
					end
				end
				else	//mux2: load input from combinational logic
				begin	
					for (x = 1; x < 10; x = x+1)
					begin
						arr[(i-1)*10 + x] <= temp[(i-1)*9 + x];	//for each cell, bits 9:1 from the combinational logic
					end
				
					if (|{&{!temp[(i-1)*9 + 1], !temp[(i-1)*9 + 2], !temp[(i-1)*9 + 3], !temp[(i-1)*9 + 4], !temp[(i-1)*9 + 5], !temp[(i-1)*9 + 6], !temp[(i-1)*9 + 7], !temp[(i-1)*9 + 8], temp[(i-1)*9 + 9]}, 
						  &{!temp[(i-1)*9 + 1], !temp[(i-1)*9 + 2], !temp[(i-1)*9 + 3], !temp[(i-1)*9 + 4], !temp[(i-1)*9 + 5], !temp[(i-1)*9 + 6], !temp[(i-1)*9 + 7], temp[(i-1)*9 + 8], !temp[(i-1)*9 + 9]},
						  &{!temp[(i-1)*9 + 1], !temp[(i-1)*9 + 2], !temp[(i-1)*9 + 3], !temp[(i-1)*9 + 4], !temp[(i-1)*9 + 5], !temp[(i-1)*9 + 6], temp[(i-1)*9 + 7], !temp[(i-1)*9 + 8], !temp[(i-1)*9 + 9]}, 
						  &{!temp[(i-1)*9 + 1], !temp[(i-1)*9 + 2], !temp[(i-1)*9 + 3], !temp[(i-1)*9 + 4], !temp[(i-1)*9 + 5], temp[(i-1)*9 + 6], !temp[(i-1)*9 + 7], !temp[(i-1)*9 + 8], !temp[(i-1)*9 + 9]}, 
						  &{!temp[(i-1)*9 + 1], !temp[(i-1)*9 + 2], !temp[(i-1)*9 + 3], !temp[(i-1)*9 + 4], temp[(i-1)*9 + 5], !temp[(i-1)*9 + 6], !temp[(i-1)*9 + 7], !temp[(i-1)*9 + 8], !temp[(i-1)*9 + 9]}, 
						  &{!temp[(i-1)*9 + 1], !temp[(i-1)*9 + 2], !temp[(i-1)*9 + 3], temp[(i-1)*9 + 4], !temp[(i-1)*9 + 5], !temp[(i-1)*9 + 6], !temp[(i-1)*9 + 7], !temp[(i-1)*9 + 8], !temp[(i-1)*9 + 9]}, 
						  &{!temp[(i-1)*9 + 1], !temp[(i-1)*9 + 2], temp[(i-1)*9 + 3], !temp[(i-1)*9 + 4], !temp[(i-1)*9 + 5], !temp[(i-1)*9 + 6], !temp[(i-1)*9 + 7], !temp[(i-1)*9 + 8], !temp[(i-1)*9 + 9]}, 
						  &{!temp[(i-1)*9 + 1], temp[(i-1)*9 + 2], !temp[(i-1)*9 + 3], !temp[(i-1)*9 + 4], !temp[(i-1)*9 + 5], !temp[(i-1)*9 + 6], !temp[(i-1)*9 + 7], !temp[(i-1)*9 + 8], !temp[(i-1)*9 + 9]}, 
						  &{temp[(i-1)*9 + 1], !temp[(i-1)*9 + 2], !temp[(i-1)*9 + 3], !temp[(i-1)*9 + 4], !temp[(i-1)*9 + 5], !temp[(i-1)*9 + 6], !temp[(i-1)*9 + 7], !temp[(i-1)*9 + 8], !temp[(i-1)*9 + 9]}})
					begin
						arr[(i-1)*10 + 10] <= 1;	//mux3: 10th bit of each cell- if one of the combinations above- set
					end
					else
					begin
						arr[(i-1)*10 + 10] <= 0;	//mux3: 10th bit of each cell- if more that one bit set, then not confirmed
					end
				end //else load
			end	//for
	end	//always @
	
	
	
endmodule



		
